//
// bootrom
//


`include "define.vh"

module bootrom (
    input wire clk,
    input wire [31:0] addr,
    output wire [31:0] rd_data
);

    //reg [31:0] mem [0:1023];  // 4KiB(12bitアドレス空間)
    wire [31:0] mem [0:638];  // 4KiB(12bitアドレス空間)
    reg [9:0] addr_sync;  // 4KiBを表現するための10bitアドレス(下位2bitはここでは考慮しない)

    //initial $readmemh({`BOOTROM_DATA_PATH, "code.hex"}, mem);

    assign mem[0] = 32'h0080006f;
    assign mem[1] = 32'h0000006f;
    assign mem[2] = 32'h00000093;
    assign mem[3] = 32'h00000113;
    assign mem[4] = 32'h00000193;
    assign mem[5] = 32'h00000213;
    assign mem[6] = 32'h00000293;
    assign mem[7] = 32'h00000313;
    assign mem[8] = 32'h00000393;
    assign mem[9] = 32'h00000413;
    assign mem[10] = 32'h00000493;
    assign mem[11] = 32'h00000513;
    assign mem[12] = 32'h00000593;
    assign mem[13] = 32'h00000613;
    assign mem[14] = 32'h00000693;
    assign mem[15] = 32'h00000713;
    assign mem[16] = 32'h00000793;
    assign mem[17] = 32'h00000813;
    assign mem[18] = 32'h00000893;
    assign mem[19] = 32'h00000913;
    assign mem[20] = 32'h00000993;
    assign mem[21] = 32'h00000a13;
    assign mem[22] = 32'h00000a93;
    assign mem[23] = 32'h00000b13;
    assign mem[24] = 32'h00000b93;
    assign mem[25] = 32'h00000c13;
    assign mem[26] = 32'h00000c93;
    assign mem[27] = 32'h00000d13;
    assign mem[28] = 32'h00000d93;
    assign mem[29] = 32'h00000e13;
    assign mem[30] = 32'h00000e93;
    assign mem[31] = 32'h00000f13;
    assign mem[32] = 32'h00000f93;
    assign mem[33] = 32'h00002137;
    assign mem[34] = 32'h20010113;
    assign mem[35] = 32'h031000ef;
    assign mem[36] = 32'hf75ff06f;
    assign mem[37] = 32'h00100793;
    assign mem[38] = 32'h02f58263;
    assign mem[39] = 32'h00059e63;
    assign mem[40] = 32'h00020737;
    assign mem[41] = 32'h05072583;
    assign mem[42] = 32'h00a797b3;
    assign mem[43] = 32'hfff7c793;
    assign mem[44] = 32'h00b7f7b3;
    assign mem[45] = 32'h04f72823;
    assign mem[46] = 32'h00008067;
    assign mem[47] = 32'h000207b7;
    assign mem[48] = 32'h0507a703;
    assign mem[49] = 32'h00a595b3;
    assign mem[50] = 32'h00e5e5b3;
    assign mem[51] = 32'h04b7a823;
    assign mem[52] = 32'h00008067;
    assign mem[53] = 32'h000207b7;
    assign mem[54] = 32'h0407a783;
    assign mem[55] = 32'h00a7d533;
    assign mem[56] = 32'h00157513;
    assign mem[57] = 32'h00008067;
    assign mem[58] = 32'h000207b7;
    assign mem[59] = 32'h0207a783;
    assign mem[60] = 32'h00100513;
    assign mem[61] = 32'h40f50533;
    assign mem[62] = 32'h00008067;
    assign mem[63] = 32'h000207b7;
    assign mem[64] = 32'h00100613;
    assign mem[65] = 32'h0207a703;
    assign mem[66] = 32'hfec70ee3;
    assign mem[67] = 32'h02a7a023;
    assign mem[68] = 32'h00008067;
    assign mem[69] = 32'h000207b7;
    assign mem[70] = 32'h0307a503;
    assign mem[71] = 32'h00855513;
    assign mem[72] = 32'h00157513;
    assign mem[73] = 32'h00008067;
    assign mem[74] = 32'h00020737;
    assign mem[75] = 32'h03072783;
    assign mem[76] = 32'h1007f793;
    assign mem[77] = 32'hfe078ce3;
    assign mem[78] = 32'h03072503;
    assign mem[79] = 32'h00100793;
    assign mem[80] = 32'h02f72823;
    assign mem[81] = 32'h0ff57513;
    assign mem[82] = 32'h00008067;
    assign mem[83] = 32'h000207b7;
    assign mem[84] = 32'h0107a703;
    assign mem[85] = 32'h04050263;
    assign mem[86] = 32'h0000b5b7;
    assign mem[87] = 32'hfc758613;
    assign mem[88] = 32'h000206b7;
    assign mem[89] = 32'hfc858593;
    assign mem[90] = 32'h0106a783;
    assign mem[91] = 32'h40e787b3;
    assign mem[92] = 32'h00f67c63;
    assign mem[93] = 32'h0106a783;
    assign mem[94] = 32'h00b70733;
    assign mem[95] = 32'hfff50513;
    assign mem[96] = 32'h40e787b3;
    assign mem[97] = 32'hfef668e3;
    assign mem[98] = 32'h0106a783;
    assign mem[99] = 32'h00e7f463;
    assign mem[100] = 32'h0106a703;
    assign mem[101] = 32'hfc051ae3;
    assign mem[102] = 32'h00008067;
    assign mem[103] = 32'h00060713;
    assign mem[104] = 32'h0cc05c63;
    assign mem[105] = 32'hfff60893;
    assign mem[106] = 32'h40a007b3;
    assign mem[107] = 32'h00500613;
    assign mem[108] = 32'h0ff5f593;
    assign mem[109] = 32'h0037f793;
    assign mem[110] = 32'h00088693;
    assign mem[111] = 32'h0d165663;
    assign mem[112] = 32'h0a078e63;
    assign mem[113] = 32'h00b50023;
    assign mem[114] = 32'h00100693;
    assign mem[115] = 32'h00150813;
    assign mem[116] = 32'h02d78263;
    assign mem[117] = 32'h00b500a3;
    assign mem[118] = 32'h00300693;
    assign mem[119] = 32'h00250813;
    assign mem[120] = 32'hffe70893;
    assign mem[121] = 32'h00d79863;
    assign mem[122] = 32'h00350813;
    assign mem[123] = 32'h00b50123;
    assign mem[124] = 32'hffd70893;
    assign mem[125] = 32'h00859613;
    assign mem[126] = 32'h40f70333;
    assign mem[127] = 32'h00c5e633;
    assign mem[128] = 32'h01059693;
    assign mem[129] = 32'h00d666b3;
    assign mem[130] = 32'h01859713;
    assign mem[131] = 32'h00f507b3;
    assign mem[132] = 32'hffc37613;
    assign mem[133] = 32'h00e6e733;
    assign mem[134] = 32'h00f606b3;
    assign mem[135] = 32'h00e7a023;
    assign mem[136] = 32'h00478793;
    assign mem[137] = 32'hfed79ce3;
    assign mem[138] = 32'hffc37693;
    assign mem[139] = 32'h40d88733;
    assign mem[140] = 32'h00d807b3;
    assign mem[141] = 32'h04d30263;
    assign mem[142] = 32'hfff70693;
    assign mem[143] = 32'h00b78023;
    assign mem[144] = 32'h02068c63;
    assign mem[145] = 32'h00b780a3;
    assign mem[146] = 32'hffe70693;
    assign mem[147] = 32'h02068663;
    assign mem[148] = 32'h00b78123;
    assign mem[149] = 32'hffd70693;
    assign mem[150] = 32'h02068063;
    assign mem[151] = 32'h00b781a3;
    assign mem[152] = 32'hffc70693;
    assign mem[153] = 32'h00068a63;
    assign mem[154] = 32'h00b78223;
    assign mem[155] = 32'h00500693;
    assign mem[156] = 32'h00d70463;
    assign mem[157] = 32'h00b782a3;
    assign mem[158] = 32'h00008067;
    assign mem[159] = 32'h00050813;
    assign mem[160] = 32'h00070893;
    assign mem[161] = 32'hf71ff06f;
    assign mem[162] = 32'h00050793;
    assign mem[163] = 32'hfb1ff06f;
    assign mem[164] = 32'h0ac05a63;
    assign mem[165] = 32'h00158693;
    assign mem[166] = 32'h40d507b3;
    assign mem[167] = 32'hfff60713;
    assign mem[168] = 32'h0037b793;
    assign mem[169] = 32'h00973713;
    assign mem[170] = 32'h0017c793;
    assign mem[171] = 32'h00174713;
    assign mem[172] = 32'h00e7f7b3;
    assign mem[173] = 32'h06078a63;
    assign mem[174] = 32'h00a5e7b3;
    assign mem[175] = 32'h0037f793;
    assign mem[176] = 32'h06079463;
    assign mem[177] = 32'hffc67813;
    assign mem[178] = 32'h00058793;
    assign mem[179] = 32'h00050713;
    assign mem[180] = 32'h00b80833;
    assign mem[181] = 32'h0007a683;
    assign mem[182] = 32'h00478793;
    assign mem[183] = 32'h00470713;
    assign mem[184] = 32'hfed72e23;
    assign mem[185] = 32'hff0798e3;
    assign mem[186] = 32'hffc67793;
    assign mem[187] = 32'h00367693;
    assign mem[188] = 32'h00f50733;
    assign mem[189] = 32'h00f585b3;
    assign mem[190] = 32'h04f60663;
    assign mem[191] = 32'h0005c603;
    assign mem[192] = 32'hfff68793;
    assign mem[193] = 32'h00c70023;
    assign mem[194] = 32'h02078e63;
    assign mem[195] = 32'h0015c603;
    assign mem[196] = 32'h00200793;
    assign mem[197] = 32'h00c700a3;
    assign mem[198] = 32'h02f68663;
    assign mem[199] = 32'h0025c783;
    assign mem[200] = 32'h00f70123;
    assign mem[201] = 32'h00008067;
    assign mem[202] = 32'h00c50633;
    assign mem[203] = 32'h00050793;
    assign mem[204] = 32'hfff6c703;
    assign mem[205] = 32'h00178793;
    assign mem[206] = 32'h00168693;
    assign mem[207] = 32'hfee78fa3;
    assign mem[208] = 32'hfec798e3;
    assign mem[209] = 32'h00008067;
    assign mem[210] = 32'h02c05a63;
    assign mem[211] = 32'h00c58633;
    assign mem[212] = 32'h0080006f;
    assign mem[213] = 32'h02b60463;
    assign mem[214] = 32'h00054783;
    assign mem[215] = 32'h0005c703;
    assign mem[216] = 32'h00150513;
    assign mem[217] = 32'h00158593;
    assign mem[218] = 32'hfee786e3;
    assign mem[219] = 32'h00f737b3;
    assign mem[220] = 32'h00179513;
    assign mem[221] = 32'hfff50513;
    assign mem[222] = 32'h00008067;
    assign mem[223] = 32'h00000513;
    assign mem[224] = 32'h00008067;
    assign mem[225] = 32'h00054783;
    assign mem[226] = 32'h00050713;
    assign mem[227] = 32'h00000513;
    assign mem[228] = 32'h00078c63;
    assign mem[229] = 32'h00150513;
    assign mem[230] = 32'h00a707b3;
    assign mem[231] = 32'h0007c783;
    assign mem[232] = 32'hfe079ae3;
    assign mem[233] = 32'h00008067;
    assign mem[234] = 32'h00008067;
    assign mem[235] = 32'h0005c703;
    assign mem[236] = 32'h00050793;
    assign mem[237] = 32'h00e50023;
    assign mem[238] = 32'h00070c63;
    assign mem[239] = 32'h0015c703;
    assign mem[240] = 32'h00178793;
    assign mem[241] = 32'h00158593;
    assign mem[242] = 32'h00e78023;
    assign mem[243] = 32'hfe0718e3;
    assign mem[244] = 32'h00008067;
    assign mem[245] = 32'h0080006f;
    assign mem[246] = 32'h02e79263;
    assign mem[247] = 32'h00054783;
    assign mem[248] = 32'h0005c703;
    assign mem[249] = 32'h00150513;
    assign mem[250] = 32'h00158593;
    assign mem[251] = 32'h00e7e6b3;
    assign mem[252] = 32'hfe0694e3;
    assign mem[253] = 32'h00000513;
    assign mem[254] = 32'h00008067;
    assign mem[255] = 32'h00f737b3;
    assign mem[256] = 32'h00179513;
    assign mem[257] = 32'hfff50513;
    assign mem[258] = 32'h00008067;
    assign mem[259] = 32'h00c50633;
    assign mem[260] = 32'h00054783;
    assign mem[261] = 32'h40a60733;
    assign mem[262] = 32'h00150513;
    assign mem[263] = 32'h00079663;
    assign mem[264] = 32'h0005c683;
    assign mem[265] = 32'h02068263;
    assign mem[266] = 32'h02e05063;
    assign mem[267] = 32'h0005c703;
    assign mem[268] = 32'h00158593;
    assign mem[269] = 32'hfcf70ee3;
    assign mem[270] = 32'h00f737b3;
    assign mem[271] = 32'h00179513;
    assign mem[272] = 32'hfff50513;
    assign mem[273] = 32'h00008067;
    assign mem[274] = 32'h00000513;
    assign mem[275] = 32'h00008067;
    assign mem[276] = 32'hff010113;
    assign mem[277] = 32'h00812423;
    assign mem[278] = 32'h00112623;
    assign mem[279] = 32'h00a00793;
    assign mem[280] = 32'h00050413;
    assign mem[281] = 32'h02f50063;
    assign mem[282] = 32'h00040513;
    assign mem[283] = 32'hc91ff0ef;
    assign mem[284] = 32'h00c12083;
    assign mem[285] = 32'h00812403;
    assign mem[286] = 32'h00000513;
    assign mem[287] = 32'h01010113;
    assign mem[288] = 32'h00008067;
    assign mem[289] = 32'h00d00513;
    assign mem[290] = 32'hc75ff0ef;
    assign mem[291] = 32'h00040513;
    assign mem[292] = 32'hc6dff0ef;
    assign mem[293] = 32'h00c12083;
    assign mem[294] = 32'h00812403;
    assign mem[295] = 32'h00000513;
    assign mem[296] = 32'h01010113;
    assign mem[297] = 32'h00008067;
    assign mem[298] = 32'hff010113;
    assign mem[299] = 32'h00812423;
    assign mem[300] = 32'h00112623;
    assign mem[301] = 32'h00912223;
    assign mem[302] = 32'h00050413;
    assign mem[303] = 32'h00054503;
    assign mem[304] = 32'h00050e63;
    assign mem[305] = 32'h00a00493;
    assign mem[306] = 32'h00140413;
    assign mem[307] = 32'h02950463;
    assign mem[308] = 32'hc2dff0ef;
    assign mem[309] = 32'h00044503;
    assign mem[310] = 32'hfe0518e3;
    assign mem[311] = 32'h00c12083;
    assign mem[312] = 32'h00812403;
    assign mem[313] = 32'h00412483;
    assign mem[314] = 32'h00000513;
    assign mem[315] = 32'h01010113;
    assign mem[316] = 32'h00008067;
    assign mem[317] = 32'h00d00513;
    assign mem[318] = 32'hc05ff0ef;
    assign mem[319] = 32'h00a00513;
    assign mem[320] = 32'hbfdff0ef;
    assign mem[321] = 32'h00044503;
    assign mem[322] = 32'hfc0510e3;
    assign mem[323] = 32'h00c12083;
    assign mem[324] = 32'h00812403;
    assign mem[325] = 32'h00412483;
    assign mem[326] = 32'h00000513;
    assign mem[327] = 32'h01010113;
    assign mem[328] = 32'h00008067;
    assign mem[329] = 32'hfe010113;
    assign mem[330] = 32'h00112e23;
    assign mem[331] = 32'h00812c23;
    assign mem[332] = 32'h00912a23;
    assign mem[333] = 32'h00010623;
    assign mem[334] = 32'h04051863;
    assign mem[335] = 32'h00059463;
    assign mem[336] = 32'h00100593;
    assign mem[337] = 32'h00b10793;
    assign mem[338] = 32'h03000713;
    assign mem[339] = 32'h00058a63;
    assign mem[340] = 32'h00e78023;
    assign mem[341] = 32'hfff58593;
    assign mem[342] = 32'hfff78793;
    assign mem[343] = 32'hfe059ae3;
    assign mem[344] = 32'h0017c503;
    assign mem[345] = 32'h00178413;
    assign mem[346] = 32'h00a00493;
    assign mem[347] = 32'h08051463;
    assign mem[348] = 32'h01c12083;
    assign mem[349] = 32'h01812403;
    assign mem[350] = 32'h01412483;
    assign mem[351] = 32'h00000513;
    assign mem[352] = 32'h02010113;
    assign mem[353] = 32'h00008067;
    assign mem[354] = 32'h00050713;
    assign mem[355] = 32'h00001837;
    assign mem[356] = 32'h00f77793;
    assign mem[357] = 32'h10c80813;
    assign mem[358] = 32'h00f807b3;
    assign mem[359] = 32'h0007c503;
    assign mem[360] = 32'h00b10413;
    assign mem[361] = 32'hfff40793;
    assign mem[362] = 32'h00a780a3;
    assign mem[363] = 32'h00475713;
    assign mem[364] = 32'h02058663;
    assign mem[365] = 32'hfff58593;
    assign mem[366] = 32'hf80708e3;
    assign mem[367] = 32'h00078413;
    assign mem[368] = 32'h00f77793;
    assign mem[369] = 32'h00f807b3;
    assign mem[370] = 32'h0007c503;
    assign mem[371] = 32'h00475713;
    assign mem[372] = 32'hfff40793;
    assign mem[373] = 32'h00a780a3;
    assign mem[374] = 32'hfc059ee3;
    assign mem[375] = 32'h00f77693;
    assign mem[376] = 32'h00d806b3;
    assign mem[377] = 32'hfff78613;
    assign mem[378] = 32'h04071c63;
    assign mem[379] = 32'h00a00493;
    assign mem[380] = 32'hf80500e3;
    assign mem[381] = 32'h00140413;
    assign mem[382] = 32'h00950c63;
    assign mem[383] = 32'hb01ff0ef;
    assign mem[384] = 32'h00044503;
    assign mem[385] = 32'hf60506e3;
    assign mem[386] = 32'h00140413;
    assign mem[387] = 32'hfe9518e3;
    assign mem[388] = 32'h00d00513;
    assign mem[389] = 32'hae9ff0ef;
    assign mem[390] = 32'h00a00513;
    assign mem[391] = 32'hae1ff0ef;
    assign mem[392] = 32'h00044503;
    assign mem[393] = 32'hfc0518e3;
    assign mem[394] = 32'h01c12083;
    assign mem[395] = 32'h01812403;
    assign mem[396] = 32'h01412483;
    assign mem[397] = 32'h00000513;
    assign mem[398] = 32'h02010113;
    assign mem[399] = 32'h00008067;
    assign mem[400] = 32'h0006c503;
    assign mem[401] = 32'h00078413;
    assign mem[402] = 32'h00475713;
    assign mem[403] = 32'h00a78023;
    assign mem[404] = 32'h00060793;
    assign mem[405] = 32'hf89ff06f;
    assign mem[406] = 32'hff010113;
    assign mem[407] = 32'h00112623;
    assign mem[408] = 32'h00812423;
    assign mem[409] = 32'hac5ff0ef;
    assign mem[410] = 32'h00d00793;
    assign mem[411] = 32'h02f50663;
    assign mem[412] = 32'h00a00793;
    assign mem[413] = 32'h00050413;
    assign mem[414] = 32'h02f50063;
    assign mem[415] = 32'h00040513;
    assign mem[416] = 32'ha7dff0ef;
    assign mem[417] = 32'h00c12083;
    assign mem[418] = 32'h00040513;
    assign mem[419] = 32'h00812403;
    assign mem[420] = 32'h01010113;
    assign mem[421] = 32'h00008067;
    assign mem[422] = 32'h00d00513;
    assign mem[423] = 32'ha61ff0ef;
    assign mem[424] = 32'h00a00413;
    assign mem[425] = 32'h00040513;
    assign mem[426] = 32'ha55ff0ef;
    assign mem[427] = 32'h00c12083;
    assign mem[428] = 32'h00040513;
    assign mem[429] = 32'h00812403;
    assign mem[430] = 32'h01010113;
    assign mem[431] = 32'h00008067;
    assign mem[432] = 32'hfe010113;
    assign mem[433] = 32'h00812c23;
    assign mem[434] = 32'h00912a23;
    assign mem[435] = 32'h01212823;
    assign mem[436] = 32'h01312623;
    assign mem[437] = 32'h01412423;
    assign mem[438] = 32'h00112e23;
    assign mem[439] = 32'h00050493;
    assign mem[440] = 32'h00d00993;
    assign mem[441] = 32'ha45ff0ef;
    assign mem[442] = 32'h00000913;
    assign mem[443] = 32'h00a00a13;
    assign mem[444] = 32'h00050413;
    assign mem[445] = 32'h03350663;
    assign mem[446] = 32'h03450463;
    assign mem[447] = 32'ha01ff0ef;
    assign mem[448] = 32'h00848023;
    assign mem[449] = 32'h00190793;
    assign mem[450] = 32'h00148493;
    assign mem[451] = 32'h02040463;
    assign mem[452] = 32'h00078913;
    assign mem[453] = 32'ha15ff0ef;
    assign mem[454] = 32'h00050413;
    assign mem[455] = 32'hfd351ee3;
    assign mem[456] = 32'h00d00513;
    assign mem[457] = 32'h9d9ff0ef;
    assign mem[458] = 32'h00a00513;
    assign mem[459] = 32'h9d1ff0ef;
    assign mem[460] = 32'h00048023;
    assign mem[461] = 32'h01c12083;
    assign mem[462] = 32'h01812403;
    assign mem[463] = 32'h01412483;
    assign mem[464] = 32'h00c12983;
    assign mem[465] = 32'h00812a03;
    assign mem[466] = 32'h00090513;
    assign mem[467] = 32'h01012903;
    assign mem[468] = 32'h02010113;
    assign mem[469] = 32'h00008067;
    assign mem[470] = 32'hfc010113;
    assign mem[471] = 32'h02912a23;
    assign mem[472] = 32'h03212823;
    assign mem[473] = 32'h03312623;
    assign mem[474] = 32'h03412423;
    assign mem[475] = 32'h03512223;
    assign mem[476] = 32'h03612023;
    assign mem[477] = 32'h01712e23;
    assign mem[478] = 32'h01812c23;
    assign mem[479] = 32'h01912a23;
    assign mem[480] = 32'h02112e23;
    assign mem[481] = 32'h02812c23;
    assign mem[482] = 32'h01a12823;
    assign mem[483] = 32'h01b12623;
    assign mem[484] = 32'h00050b13;
    assign mem[485] = 32'h00100993;
    assign mem[486] = 32'h00000b93;
    assign mem[487] = 32'h00000493;
    assign mem[488] = 32'h00018c37;
    assign mem[489] = 32'h00400913;
    assign mem[490] = 32'h01800a13;
    assign mem[491] = 32'h00100a93;
    assign mem[492] = 32'h0ff00c93;
    assign mem[493] = 32'h00048c63;
    assign mem[494] = 32'h971ff0ef;
    assign mem[495] = 32'h03250a63;
    assign mem[496] = 32'h03450e63;
    assign mem[497] = 32'h07550e63;
    assign mem[498] = 32'h02049a63;
    assign mem[499] = 32'h6a0c0413;
    assign mem[500] = 32'h0080006f;
    assign mem[501] = 32'h0c040e63;
    assign mem[502] = 32'h93dff0ef;
    assign mem[503] = 32'hfff40413;
    assign mem[504] = 32'hfe050ae3;
    assign mem[505] = 32'h00000493;
    assign mem[506] = 32'h941ff0ef;
    assign mem[507] = 32'hfd251ae3;
    assign mem[508] = 32'h00600513;
    assign mem[509] = 32'h909ff0ef;
    assign mem[510] = 32'h0080006f;
    assign mem[511] = 32'hfff00b93;
    assign mem[512] = 32'h03c12083;
    assign mem[513] = 32'h03812403;
    assign mem[514] = 32'h03412483;
    assign mem[515] = 32'h03012903;
    assign mem[516] = 32'h02c12983;
    assign mem[517] = 32'h02812a03;
    assign mem[518] = 32'h02412a83;
    assign mem[519] = 32'h02012b03;
    assign mem[520] = 32'h01812c03;
    assign mem[521] = 32'h01412c83;
    assign mem[522] = 32'h01012d03;
    assign mem[523] = 32'h00c12d83;
    assign mem[524] = 32'h000b8513;
    assign mem[525] = 32'h01c12b83;
    assign mem[526] = 32'h04010113;
    assign mem[527] = 32'h00008067;
    assign mem[528] = 32'h8e9ff0ef;
    assign mem[529] = 32'h00148493;
    assign mem[530] = 32'h05351e63;
    assign mem[531] = 32'h8ddff0ef;
    assign mem[532] = 32'h013547b3;
    assign mem[533] = 32'h0ff7f793;
    assign mem[534] = 32'h05979663;
    assign mem[535] = 32'h080b0413;
    assign mem[536] = 32'h000b0d93;
    assign mem[537] = 32'h00000d13;
    assign mem[538] = 32'h8c1ff0ef;
    assign mem[539] = 32'h001d8d93;
    assign mem[540] = 32'h01a50d33;
    assign mem[541] = 32'hfead8fa3;
    assign mem[542] = 32'h0ffd7d13;
    assign mem[543] = 32'hffb416e3;
    assign mem[544] = 32'h8a9ff0ef;
    assign mem[545] = 32'h02ad1063;
    assign mem[546] = 32'h00198993;
    assign mem[547] = 32'h00600513;
    assign mem[548] = 32'h0ff9f993;
    assign mem[549] = 32'h080b8b93;
    assign mem[550] = 32'h865ff0ef;
    assign mem[551] = 32'h00040b13;
    assign mem[552] = 32'hf15ff06f;
    assign mem[553] = 32'h01500513;
    assign mem[554] = 32'h855ff0ef;
    assign mem[555] = 32'hf09ff06f;
    assign mem[556] = 32'h01500513;
    assign mem[557] = 32'h849ff0ef;
    assign mem[558] = 32'hf15ff06f;
    assign mem[559] = 32'hfc010113;
    assign mem[560] = 32'h02812c23;
    assign mem[561] = 32'h02912a23;
    assign mem[562] = 32'h03212823;
    assign mem[563] = 32'h03312623;
    assign mem[564] = 32'h03412423;
    assign mem[565] = 32'h03512223;
    assign mem[566] = 32'h03612023;
    assign mem[567] = 32'h01712e23;
    assign mem[568] = 32'h01812c23;
    assign mem[569] = 32'h01912a23;
    assign mem[570] = 32'h01a12823;
    assign mem[571] = 32'h01b12623;
    assign mem[572] = 32'h02112e23;
    assign mem[573] = 32'h000019b7;
    assign mem[574] = 32'h00002437;
    assign mem[575] = 32'h00001937;
    assign mem[576] = 32'h000014b7;
    assign mem[577] = 32'h00001a37;
    assign mem[578] = 32'h00001bb7;
    assign mem[579] = 32'h00001b37;
    assign mem[580] = 32'h00001cb7;
    assign mem[581] = 32'h00001ab7;
    assign mem[582] = 32'h00001c37;
    assign mem[583] = 32'h00001db7;
    assign mem[584] = 32'h00001d37;
    assign mem[585] = 32'h00098513;
    assign mem[586] = 32'hb81ff0ef;
    assign mem[587] = 32'ha0040513;
    assign mem[588] = 32'hd91ff0ef;
    assign mem[589] = 32'h00890593;
    assign mem[590] = 32'ha0040513;
    assign mem[591] = 32'ha99ff0ef;
    assign mem[592] = 32'h00050793;
    assign mem[593] = 32'h20048513;
    assign mem[594] = 32'h00079e63;
    assign mem[595] = 32'he0dff0ef;
    assign mem[596] = 32'h00050793;
    assign mem[597] = 32'h010a0513;
    assign mem[598] = 32'h0207dc63;
    assign mem[599] = 32'hb4dff0ef;
    assign mem[600] = 32'hfc5ff06f;
    assign mem[601] = 32'h048b0593;
    assign mem[602] = 32'ha0040513;
    assign mem[603] = 32'ha69ff0ef;
    assign mem[604] = 32'h00050793;
    assign mem[605] = 32'h054a8593;
    assign mem[606] = 32'ha0040513;
    assign mem[607] = 32'h02079063;
    assign mem[608] = 32'h04cc8513;
    assign mem[609] = 32'hb25ff0ef;
    assign mem[610] = 32'h079000ef;
    assign mem[611] = 32'hf99ff06f;
    assign mem[612] = 32'h02cb8513;
    assign mem[613] = 32'hb15ff0ef;
    assign mem[614] = 32'hf8dff06f;
    assign mem[615] = 32'ha39ff0ef;
    assign mem[616] = 32'h00050793;
    assign mem[617] = 32'h060c0513;
    assign mem[618] = 32'h04079263;
    assign mem[619] = 32'hafdff0ef;
    assign mem[620] = 32'h07cd8513;
    assign mem[621] = 32'haf5ff0ef;
    assign mem[622] = 32'h094d0513;
    assign mem[623] = 32'haedff0ef;
    assign mem[624] = 32'h094d0513;
    assign mem[625] = 32'hae5ff0ef;
    assign mem[626] = 32'h000017b7;
    assign mem[627] = 32'h0ac78513;
    assign mem[628] = 32'had9ff0ef;
    assign mem[629] = 32'h000017b7;
    assign mem[630] = 32'h0c878513;
    assign mem[631] = 32'hacdff0ef;
    assign mem[632] = 32'h000017b7;
    assign mem[633] = 32'h0e478513;
    assign mem[634] = 32'hf75ff06f;
    assign mem[635] = 32'h000017b7;
    assign mem[636] = 32'h10078513;
    assign mem[637] = 32'hab5ff0ef;
    assign mem[638] = 32'hf2dff06f;
     
    always @(posedge clk) begin
        addr_sync <= addr[11:2];  // 読み出しアドレス更新をクロックと同期することでBRAM化
    end
    
    assign rd_data = mem[addr_sync];

endmodule
